module oneshot_universal(clk, rst, btn, btn_trig);
parameter WIDTH=1;
input clk, rst;
input [WIDTH-1:0] btn;
output reg [WIDTH-1:0] btn_trig;
reg [WIDTH-1:0] btn_reg;

always @(negedge rst or posedge clk) begin
    if(!rst) begin
        btn_reg <= {WIDTH{1'b0}};
        btn_trig <= {WIDTH{1'b0}};
    end else begin
        btn_reg <= btn;
        btn_trig <= btn & ~btn_reg;
    end
end
endmodule
